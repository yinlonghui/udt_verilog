﻿module	ACKtimer_top ;







endmodule