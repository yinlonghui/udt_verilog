﻿module	ProcessACK_top ;






endmodule