﻿//%	@file	CacheManager.v
//%	@brief	本文定义缓存管理

//%	
//%	@details

module CacheManager(
	input	core_clk,									//%	核心模块时钟
	input	core_rst_n,									//%	核心模块复位(低信号复位)
);



endmodule