﻿module	connect;


endmodule