﻿module	ProcessNAK_top ; 







endmodule