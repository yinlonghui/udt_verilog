﻿module SND_top ;

endmodule