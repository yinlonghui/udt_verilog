﻿//%	@file	NACKtimer.v
//%	@brief	本文件定义NACKtimer模块

//%	NACKtimer模块是NACK包计数器


module	NACKtimer(

);




endmodule