﻿//%	@file	EXPtimer.v
//%	@brief	本文件定义EXPtimer模块

//%	NACKtimer模块是EXP包计数器


module	EXPtimer(
	input	core_clk	,	//%	时钟信号
	input	core_rst_n	,	//%	时钟复位信号(低有效)

);




endmodule