﻿//%	@file	Arbitrator.v
//%	@brief	本文件定义Arbitrator模块

//%	Arbitrator 模块是ACK包计数器

module	Arbitrator(
	input	core_clk	,	//%	时钟信号
	input	core_rst_n	,	//%	时钟复位信号(低有效)

);



endmodule