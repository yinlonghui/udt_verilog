﻿module	RcvBufferManager_top ;




endmodule