﻿module  close_top ;


endmodule