﻿module	ProcessACK2_top ;






endmodule