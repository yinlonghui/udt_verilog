﻿module cc_top;





endmodule