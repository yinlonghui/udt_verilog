module	StateManager_top ;



endmodule