﻿module	decode_top;



endmodule

