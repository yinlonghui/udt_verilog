﻿module	EXPtimer_top ;




endmodule