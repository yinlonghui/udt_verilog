﻿module	mutexValue_top ;


endmodule