﻿module	SocketManager_top ;

endmodule