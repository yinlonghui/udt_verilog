﻿module	Arbitrator_top;



endmodule