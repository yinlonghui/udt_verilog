﻿//%	@file	bufferManager.v
//%	@brief	本文件定义bufferManager模块

//%	@brief	PktTimeWindow模块用于管理PktTimeWindow

module	ACKWindows(
	input	core_clk	,	//%	时钟信号
	input	core_rst_n	,	//%	时钟复位信号(低有效)

);



endmodule