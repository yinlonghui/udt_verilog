﻿//% @file   configure.v
//%	@brief	 本文件定义配置寄存器模块
//% @details 


//% 配置寄存器模块主要接收用户配置命令，以AXI-LITE协议操作BRAM，用户通过操作UDT寄存器来管理UDT
//% @details
//%	配置参数：
//%		1、配置状态寄存器标识为成功再进行2步骤
//%		2、检查是否已经UDT建立连接:
//%			2.1若已经建立连接，则将配置状态寄存器表示错误状态（连接）
//%			2.2 若未建立连接，则检查参数是否在正确的范围内
//%				2.2.1 若在正确的范围，则向写入相应的参数，然后将配置状态寄存器标识为成功配置
//%				2.2.2 若不在正确的范围，则将配置状态寄存器表示错误状态（越界）
//%	建立连接:
//%		检查连接寄存器的状态：
//%			1、若UDT连接状态寄存器为正在连接或者连接成功状态，则将UDT连接状态寄存器改为连接失败，发送给Socket Manager关闭连接的操作
//%			2、若UDT连接状态寄存器为关闭状态或者未打开状态，将UDT连接状态寄存器改为正在连接状态，发送给Socket Manager打开连接的操作
//%	关闭连接：
//%			1、若UDT连接状态为关闭，则将UDT连接状态寄存器改为关闭失败
//%			2、若UDT连接状态为连接，向Socket Manager发送关闭连接操作，等待UDT关闭，更新连接寄存器标识为关闭
//%	读状态寄存器：
//%			AXI-LITE（读操作）直接读取BRAM
//%	寄存器映射：
module    configure #(
		parameter	DEFAULT_SND_BUFFER_SIZE	=	8192 ,
		parameter	DEFAULT_REV_BUFFER_SIZE =   8192 ,
		parameter	DEFAULT_FLIGHT_FLAG_SIZE =	256000,
		parameter	DEFAULT_INIT_SEQ	=	0	,
		parameter	MAX_DDR3_SIZE	 =	1024*1024*1024*8 ,
		parameter	MAX_MSSize	= 8000	
)(
	input	ctrl_s_axi_aclk,							//% 用户-时钟信号
	input   ctrl_s_axi_aresetn,							//% 用户-复位信号
	input	[31:0]	ctrl_s_axi_awaddr,					//%	用户-写地址信号
	input	ctrl_s_axi_awvalid,							//% 用户-写地址有效
	output	ctrl_s_axi_awready,							//%	用户-写地址就绪
	input	[31:0]	ctrl_s_axi_wdata,					//%	用户-写操作数据
	input	[3:0]	ctrl_s_axi_wstrb,					//%	用户-写操作字节使能
	input	ctrl_s_axi_wvalid,							//%	用户-写数据有效
	output	ctrl_s_axi_wready,							//%	用户-写数据就绪
	output	[1:0]	ctrl_s_axi_bresp,					//%	用户-写数据应答
	output	ctrl_s_axi_bvalid,							//%	用户-写应答有效
	input	ctrl_s_axi_bready,							//%	用户-写应答就绪
	input   [31:0]	ctrl_s_axi_araddr,					//% 用户-读地址信号
	input	ctrl_s_axi_arvalid,							//% 用户-读地址有效
	output	ctrl_s_axi_arready,							//% 用户-读地址就绪
	output  [31:0]	ctrl_s_axi_rdata,					//%	用户-读操作数据
	output	[1:0]	ctrl_s_axi_rresp,					//%	用户-读数据应答
	output	ctrl_s_axi_rvalid,							//%	用户-读数据有效
	input	ctrl_s_axi_rready,							//%	用户-读数据就绪


	input	core_clk,									//%	核心模块时钟
	input	core_rst_n,									//%	核心模块复位(低信号复位)	
	input	[31:0]	udt_state ,							//%	连接状态
	input	state_valid,								//%	连接状态有效
	output	state_ready,								//%	连接状态就绪
	output	Req_Connect ,								//%	连接请求
	input	Res_Connect ,								//% 连接回应
	output	Req_Close	,								//%	关闭请求
	input	Res_Close	,								//%	关闭回应
	output	[31:0]	Snd_Buffer_Size ,					//%	发送buffer大小
	output	[31:0]	Rev_Buffer_Size	,					//%	接收buffer大小
	output	[31:0]	FlightFlagSize ,					//%	最大流量窗口大小
	output	[31:0]	MSSize								//%	最大包大小

);
/*			(Snd_Buffer_Size +   Snd_Buffer_Size)*MSSize +   2*m_iFlightFlagSize*sizeof(list) < DEFAULT_FLIGHT_FLAG_SIZE */



endmodule