﻿//% @file   udt.v
//% @brief  UDT模块

module  udt(
	input	clk ,//%  时钟
	input   rst ,//%  复位
);

endmodule