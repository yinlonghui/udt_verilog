﻿module	state2axis_top

endmodule