﻿//%	@file	list.v
//%	@brief	本文件定义list模块

//%	@brief	list模块用于管理丢失链表

module	list(
	input	core_clk	,	//%	时钟信号
	input	core_rst_n	,	//%	时钟复位信号(低有效)

);



endmodule