﻿module	ProcessClose_top;



endmodule