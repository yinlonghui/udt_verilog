﻿module   configure_top ;



endmodule