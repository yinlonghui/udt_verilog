﻿module ClientManager_top ;


endmodule