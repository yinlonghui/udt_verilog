﻿module ServerManager_top ;






endmodule