﻿module	RcvLossList_top ;



endmodule