﻿module ProcessData_top ;






endmodule