module	SNDtimer_top;


endmodule