﻿//%	@file	ACKWindows.v
//%	@brief	本文件定义ACKWindows模块

//%	@brief	ACKWindows模块用于管理ACKWindows

module	ACKWindows(
	input	core_clk	,	//%	时钟信号
	input	core_rst_n	,	//%	时钟复位信号(低有效)

);



endmodule