﻿module	ACKWindows_top;





endmodule