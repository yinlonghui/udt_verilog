﻿module	trans_keep_top ;

endmodule