﻿module	ProcessKeepAlive_top ;






endmodule