﻿module	SndBufferManager_top ;



endmodule