﻿module CacheManager_top;



endmodule