﻿//%	@file	ACKtimer.v
//%	@brief	本文件定义ACKtimer模块

//%	ACKtimer模块是ACK包计数器

module	ACKtimer(
	input	core_clk	,	//%	时钟信号
	input	core_rst_n	,	//%	时钟复位信号(低有效)

);



endmodule