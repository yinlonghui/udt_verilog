//%	@file	SNDtimer.v
//%	@brief	���ļ�����SNDtimerģ��

//%	SNDtimerģ����EXP��������

module	SNDtimer(
	input	core_clk	,	//%	ʱ���ź�
	input	core_rst_n	,	//%	ʱ�Ӹ�λ�ź�(����Ч)

);


endmodule