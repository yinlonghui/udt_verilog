﻿module	listen_top;



endmodule