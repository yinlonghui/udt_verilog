﻿module	SndLossList_top ;



endmodule