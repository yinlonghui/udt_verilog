﻿//%	@file	SND.v
//%	@brief	本文件定义SND模块

//%	SND模块是发送模块
module SND(
	input	core_clk	,	//%	时钟信号
	input	core_rst_n	,	//%	时钟复位信号(低有效)
	
);





endmodule