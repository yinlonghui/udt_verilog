﻿//%	@file	cc.v
//%	@brief	本文件定义CC模块

//%	@brief	CC模块为拥塞控制模块，现阶段暂时还有选定采用那种拥塞函数
module(
	input	core_clk	,	//%	时钟信号
	input	core_rst_n	,	//%	时钟复位信号(低有效)

	input	bSlowStart	,	//% 满速度
);





endmodule