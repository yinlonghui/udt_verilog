﻿module	udt_core_top ;

endmodule