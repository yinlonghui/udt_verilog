

interface	Socketif(	input	clk , output logic finish , output  logic err	)